*

.subckt Grovie

.model __Q1 NPN bf=200
.model __Q3 NPN bf=200
.model __Q2 NPN bf=200
.model __RV1 potentiometer( r=100k position=1 )
Q1 Net-_Q1-C_ Net-_Q1-B_ Net-_Q1-E_ __Q1
R4 VCC Net-_Q1-C_ 6.8k
R3 Net-_Q1-B_ Net-_C3-Pad1_ 390k
C2 Net-_C1-Pad1_ Net-_Q1-B_ 100n
R2 Net-_R1-Pad1_ Net-_C1-Pad1_ 8.2k
R1 Net-_R1-Pad1_ GND 1Meg
C1 Net-_C1-Pad1_ GND 68p
R19 VCC Net-_C3-Pad1_ 10k
R9 GND Net-_C3-Pad1_ 47k
C3 Net-_C3-Pad1_ GND 22u
C5 GND Net-_Q2-B_ 220n
R15 GND Net-_Q3-E_ 22k
Q3 VCC Net-_Q3-B_ Net-_Q3-E_ __Q3
R16 Net-_C4-Pad1_ Net-_Q3-E_ 2.7k
R5 Net-_Q1-E_ GND 75k
R7 Net-_Q2-B_ Net-_C3-Pad1_ 330k
R6 VCC Net-_Q2-C_ 6.8k
Q2 Net-_Q2-C_ Net-_Q2-B_ Net-_Q1-E_ __Q2
R8 Net-_Q1-C_ Net-_Q3-B_ 2.7k
C4 Net-_C4-Pad1_ Net-_C4-Pad2_ 2.2u
ARV1 GND Output1 Net-_C4-Pad2_ __RV1
R17 Output1 GND 20k
V1 VCC GND DC 9 
R10 Input1 Net-_R1-Pad1_ 5.6k
V2 Input1 GND DC 0 SIN( 0 150m 220 0 0 0 ) AC 1
.ends
